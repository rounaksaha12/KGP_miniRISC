`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:27:04 10/26/2022 
// Design Name: 
// Module Name:    DIFF_32bit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module DIFF_32bit(a,b,DIFFout);
input [31:0] a,b;
output [31:0] DIFFout;

/*incomplete module, passes the value of a as output*/
assign DIFFout=a;

endmodule
